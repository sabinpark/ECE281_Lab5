library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity ROM_176x4 is
  port (Clock : in std_logic;
  		CS_L : in std_logic;
        R_W  : in std_logic;
        Addr   : in std_logic_vector(7 downto 0);
        Data  : out std_logic_vector(3 downto 0));
end ROM_176x4;

architecture ROM_176x4_Arch of ROM_176x4 is
  type rom_type is array (0 to 175)
        of std_logic_vector (3 downto 0);
  signal ROM : rom_type;
  signal Read_Enable : std_logic;
begin

ROM(0) <= X"7";
ROM(1) <= X"0";
ROM(2) <= X"D";
ROM(3) <= X"2";
ROM(4) <= X"B";
ROM(5) <= X"D";
ROM(6) <= X"1";
ROM(7) <= X"B";
ROM(8) <= X"4";
ROM(9) <= X"1";
ROM(10) <= X"4";
ROM(11) <= X"2";
ROM(12) <= X"5";
ROM(13) <= X"0";
ROM(14) <= X"B";
ROM(15) <= X"E";
ROM(16) <= X"4";
ROM(17) <= X"F";
ROM(18) <= X"2";
ROM(19) <= X"B";
ROM(20) <= X"6";
ROM(21) <= X"1";
ROM(22) <= X"D";
ROM(23) <= X"2";
ROM(24) <= X"B";
ROM(25) <= X"4";
ROM(26) <= X"2";
ROM(27) <= X"6";
ROM(28) <= X"7";
ROM(29) <= X"A";
ROM(30) <= X"3";
ROM(31) <= X"2";
ROM(32) <= X"9";
ROM(33) <= X"C";
ROM(34) <= X"0";
ROM(35) <= X"F";
ROM(36) <= X"1";
ROM(37) <= X"B";
ROM(38) <= X"6";
ROM(39) <= X"7";
ROM(40) <= X"A";
ROM(41) <= X"F";
ROM(42) <= X"3";
ROM(43) <= X"7";
ROM(44) <= X"0";
ROM(45) <= X"D";
ROM(46) <= X"2";
ROM(47) <= X"B";
ROM(48) <= X"4";
ROM(49) <= X"2";
ROM(50) <= X"F";
ROM(51) <= X"1";
ROM(52) <= X"B";
ROM(53) <= X"6";
ROM(54) <= X"1";
ROM(55) <= X"D";
ROM(56) <= X"1";
ROM(57) <= X"B";
ROM(58) <= X"4";
ROM(59) <= X"1";
ROM(60) <= X"9";
ROM(61) <= X"C";
ROM(62) <= X"0";
ROM(63) <= X"7";
ROM(64) <= X"0";
ROM(65) <= X"D";
ROM(66) <= X"2";
ROM(67) <= X"B";
ROM(68) <= X"D";
ROM(69) <= X"1";
ROM(70) <= X"B";
ROM(71) <= X"4";
ROM(72) <= X"1";
ROM(73) <= X"4";
ROM(74) <= X"2";
ROM(75) <= X"9";
ROM(76) <= X"C";
ROM(77) <= X"0";
ROM(78) <= X"5";
ROM(79) <= X"0";
ROM(80) <= X"B";
ROM(81) <= X"6";
ROM(82) <= X"5";
ROM(83) <= X"9";
ROM(84) <= X"C";
ROM(85) <= X"0";
ROM(86) <= X"F";
ROM(87) <= X"2";
ROM(88) <= X"B";
ROM(89) <= X"A";
ROM(90) <= X"6";
ROM(91) <= X"6";
ROM(92) <= X"6";
ROM(93) <= X"F";
ROM(94) <= X"D";
ROM(95) <= X"2";
ROM(96) <= X"B";
ROM(97) <= X"4";
ROM(98) <= X"2";
ROM(99) <= X"9";
ROM(100) <= X"E";
ROM(101) <= X"4";
ROM(102) <= X"F";
ROM(103) <= X"1";
ROM(104) <= X"B";
ROM(105) <= X"A";
ROM(106) <= X"D";
ROM(107) <= X"7";
ROM(108) <= X"6";
ROM(109) <= X"F";
ROM(110) <= X"D";
ROM(111) <= X"1";
ROM(112) <= X"B";
ROM(113) <= X"4";
ROM(114) <= X"1";
ROM(115) <= X"7";
ROM(116) <= X"9";
ROM(117) <= X"D";
ROM(118) <= X"2";
ROM(119) <= X"B";
ROM(120) <= X"4";
ROM(121) <= X"2";
ROM(122) <= X"9";
ROM(123) <= X"E";
ROM(124) <= X"4";
ROM(125) <= X"7";
ROM(126) <= X"9";
ROM(127) <= X"D";
ROM(128) <= X"1";
ROM(129) <= X"B";
ROM(130) <= X"D";
ROM(131) <= X"2";
ROM(132) <= X"B";
ROM(133) <= X"4";
ROM(134) <= X"2";
ROM(135) <= X"4";
ROM(136) <= X"1";
ROM(137) <= X"9";
ROM(138) <= X"E";
ROM(139) <= X"4";
ROM(140) <= X"0";
ROM(141) <= X"0";
ROM(142) <= X"0";
ROM(143) <= X"0";
ROM(144) <= X"0";
ROM(145) <= X"0";
ROM(146) <= X"0";
ROM(147) <= X"0";
ROM(148) <= X"0";
ROM(149) <= X"0";
ROM(150) <= X"0";
ROM(151) <= X"0";
ROM(152) <= X"0";
ROM(153) <= X"0";
ROM(154) <= X"0";
ROM(155) <= X"0";
ROM(156) <= X"0";
ROM(157) <= X"0";
ROM(158) <= X"0";
ROM(159) <= X"0";
ROM(160) <= X"0";
ROM(161) <= X"0";
ROM(162) <= X"0";
ROM(163) <= X"0";
ROM(164) <= X"0";
ROM(165) <= X"0";
ROM(166) <= X"0";
ROM(167) <= X"0";
ROM(168) <= X"0";
ROM(169) <= X"0";
ROM(170) <= X"0";
ROM(171) <= X"0";
ROM(172) <= X"0";
ROM(173) <= X"0";
ROM(174) <= X"0";
ROM(175) <= X"0";
	Read_Enable <=  '0' when(CS_L='0' and R_W = '1') else '1';

	process (Clock)
	begin
		if(Clock='0') then
			if(Read_Enable = '0') then
			  Data  <= ROM(conv_integer(Addr));
		  	else
			  Data <= "ZZZZ";
	      	end if;
		else Data <= "ZZZZ";
		end if;

	end process;

	end ROM_176x4_Arch;
